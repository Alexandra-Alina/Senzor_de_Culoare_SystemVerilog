`ifndef TEST_PKG_SV
`define TEST_PKG_SV

package test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "test_base.sv"
  
endpackage:test_pkg

`endif