`ifndef APB_PKG_SV
`define APB_PKG_SV

package apb_pkg;

   import uvm_pkg::*;
   `include "uvm_macros.svh"

   `include "apb_defines.sv"
   `include "apb_types.sv"
   `include "apb_trans.sv"
   `include "apb_monitor.sv"
   `include "apb_sequencer.sv"
   `include "apb_seq_lib.sv"
   `include "apb_driver.sv"
   `include "apb_agent.sv"
   `include "apb_coverage.sv"
    
endpackage : apb_pkg

`endif