`define APB_AW 5
`define APB_DW 32