`ifndef APB_TYPES_SV
`define APB_TYPES_SV

typedef enum { APB_WRITE, APB_READ } apb_access_kind_t;

`endif

