`define I2C_AW 7
`define I2C_DW 8