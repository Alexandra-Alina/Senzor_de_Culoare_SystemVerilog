
  `include "test_base.sv"
  `include "test_registers.sv"
